
`ifndef __TB_PACKAGE_SV__
 `define __TB_PACKAGE_SV__
package tb_package;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "example_data_item.svh"
  `include "example_data_item2.svh"
  `include "example_seq0.svh"
  `include "example_seq1.svh"
  `include "monitor.svh"
  `include "driver.svh"
  `include "agent.svh"
  `include "scoreboard.svh"
  `include "env.svh"
endpackage: tb_package
`endif 
